CircuitMaker Text
5.6
Probes: 1
R1_1
Operating Point
0 262 142 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 10
1207 516 1913 1272
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1207 894 1913 1272
9961490 0
0
6 Title:
5 Name:
0
0
0
5
9 I Source~
198 193 71 0 2 5
0 5 4
0
0 0 17264 90
5 100mA
-18 -20 17 -12
3 Is1
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 0 0 0 0
2 Is
8157 0 0
2
44359.1 0
0
7 Ground~
168 197 232 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5572 0 0
2
44359.1 1
0
9 V Source~
197 122 142 0 2 5
0 5 2
0
0 0 17264 0
3 10V
13 0 34 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8901 0 0
2
44359.1 0
0
9 Resistor~
219 260 172 0 3 5
0 2 3 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
44359.1 0
0
9 Resistor~
219 260 97 0 2 5
0 3 4
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4747 0 0
2
44359.1 2
0
5
1 2 3 0 0 4224 0 5 4 0 0 2
260 115
260 154
1 0 2 0 0 8192 0 4 0 0 5 3
260 190
260 196
197 196
2 2 4 0 0 4224 0 1 5 0 0 3
214 71
260 71
260 79
1 1 5 0 0 4224 0 3 1 0 0 3
122 121
122 71
172 71
1 2 2 0 0 8320 0 2 3 0 0 4
197 226
197 196
122 196
122 163
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
54 259 147 283
60 263 140 279
10 this sucks
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
